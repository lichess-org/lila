playWithAFriend=Spela med en vän
inviteAFriendToPlayWithYou=Bjud in en vän att spela med dig
playWithTheMachine=Spela mot datorn
challengeTheArtificialIntelligence=Utmana datorn
toInviteSomeoneToPlayGiveThisUrl=För att bjuda in någon att spela, ge dem den här länken
gameOver=Partiet är slut
waitingForOpponent=Väntar på motståndare
waiting=Väntar
yourTurn=Din tur
aiNameLevelAiLevel=%s nivå %s
level=Nivå
toggleTheChat=Dölj/visa chattrutan
toggleSound=Ljud av/på
chat=Chatt
resign=Ge upp
checkmate=Schackmatt
stalemate=Patt
white=Vit
black=Svart
randomColor=Slumpa färg
createAGame=Skapa ett parti
whiteIsVictorious=Vit vinner
blackIsVictorious=Svart vinner
playWithTheSameOpponentAgain=Spela mot samma motståndare igen
newOpponent=Ny motståndare
playWithAnotherOpponent=Spela mot en annan motståndare
yourOpponentWantsToPlayANewGameWithYou=Din motståndare vill spela ett nytt parti med dig
joinTheGame=Starta partiet
whitePlays=Vits drag
blackPlays=Svart drag
theOtherPlayerHasLeftTheGameYouCanForceResignationOrWaitForHim=Den andre spelaren har lämnat partiet. Du kan ta en vinst, ta remi eller vänta på honom.
makeYourOpponentResign=Tvinga din motståndare att ge upp
forceResignation=Ta en vinst
forceDraw=Ta remi
talkInChat=Prata i chatten
theFirstPersonToComeOnThisUrlWillPlayWithYou=Den första som använder den här länken kommer att spela med dig
whiteCreatesTheGame=Vit startar ett parti
blackCreatesTheGame=Svart startar ett parti
whiteJoinsTheGame=Vit ansluter till partiet
blackJoinsTheGame=Svart ansluter till partiet
whiteResigned=Vit har gett upp
blackResigned=Svart har gett upp
whiteLeftTheGame=Vit har lämnat partiet
blackLeftTheGame=Svart har lämnat partiet
shareThisUrlToLetSpectatorsSeeTheGame=Dela den här länken så åskådare kan se spelet
youAreViewingThisGameAsASpectator=Du tittar på spelet som åskådare
replayAndAnalyse=Visa repris och analysera
computerAnalysisInProgress=Datorn analyserar
theComputerAnalysisYouRequestedIsNowAvailable=Datoranalysen som du begärde är nu tillgänglig
theComputerAnalysisHasFailed=Datoranalysen misslyckades
viewTheComputerAnalysis=Visa datoranalysen
requestAComputerAnalysis=Begär en datoranalys
blunders=Blunder
mistakes=Misstag
inaccuracies=Felaktighet
viewGameStats=Visa statistik
flipBoard=Vänd brädet
threefoldRepetition=Trefaldig upprepning
claimADraw=Ta remi
offerDraw=Föreslå remi
draw=Remi
nbConnectedPlayers=%s anslutna spelare
talkAboutChessAndDiscussLichessFeaturesInTheForum=Prata om schack och diskutera sidans funktioner i forumet
seeTheGamesBeingPlayedInRealTime=Se de partier som spelas i realtid
gamesBeingPlayedRightNow=Partier som spelas just nu
viewAllNbGames=Visa alla %s partier
viewNbCheckmates=Visa %s  schackmatt
nbBookmarks=%s Bokmärken
nbPopularGames=%s Populära Spel
nbAnalysedGames=%s Spelen Analyserades
bookmarkedByNbPlayers=Bokmärkt av %s spelare
viewInFullSize=Visa i full storlek
logOut=Logga ut
signIn=Logga in
newToLichess=Ny användare?
youNeedAnAccountToDoThat=Du behöver ett konto för att göra det
signUp=Registrera dig
games=Partier
forum=Forum
xPostedInForumY=%s postade i forumet %s
players=Schackspelare
minutesPerSide=Minuter per spelare
variant=Variant
timeControl=Tidskontroll
time=Tid
username=Användarnamn
password=Lösenord
haveAnAccount=Har du ett konto?
allYouNeedIsAUsernameAndAPassword=Allt du behöver är ett användarnamn och ett lösenord.
changePassword=Ändra lösenord
learnMoreAboutLichess=Lär mer om Lichess
rank=Rankning
gamesPlayed=Partier spelade
nbGamesWithYou=%s partin med dig
declineInvitation=Avböj inbjudan
cancel=Avbryt
timeOut=Time out
drawOfferSent=Remi föreslagen
drawOfferDeclined=Remi nekad
drawOfferAccepted=Remi accepterad
drawOfferCanceled=Remiförfrågan avbruten
yourOpponentOffersADraw=Din motståndare bjuder remi
accept=Acceptera
decline=Avböj
playingRightNow=Spelar nu
finished=Klart
abortGame=Avsluta parti
gameAborted=Parti avslutat
standard=Standard
unlimited=Obegränsad
mode=Läge
casual=Casual
rated=Poängsatt
thisGameIsRated=Detta parti spelas om ranking
rematch=Returmatch
rematchOfferSent=Förslag om returmatch skickat
rematchOfferAccepted=Förslag om returmatch accepterat
rematchOfferCanceled=Anbud om returmatch avbrutet
rematchOfferDeclined=Anbud om returmatch avböjt
cancelRematchOffer=Avbryt returmatchförslag
viewRematch=Visa returmatch
play=Spela
inbox=Inkorg
chatRoom=Chattrum
spectatorRoom=Åskådarrum
composeMessage=Sammanställ meddelande
noNewMessages=Inga nya meddelanden
subject=Ämne
recipient=Mottagare
send=Skicka
incrementInSeconds=Ökning i sekunder
freeOnlineChess=Gratis Schack på internet
spectators=Åskådare
nbWins=%s vinster
nbLosses=%s förluster
nbDraws=%s remi
exportGames=Exportera spel
color=Färg
ratingRange=Elo spann
giveNbSeconds=Ge  %s sekunder
premoveEnabledClickAnywhereToCancel=Premove är på -Klicka var som helst för att avbryta
thisPlayerUsesChessComputerAssistance=Den här spelaren tar hjälp av schackmotor
opening=Öppning
takeback=Bakåtsteg
proposeATakeback=Föreslå bakåtsteg
takebackPropositionSent=Förslag på bakåtsteg skickat
takebackPropositionDeclined=Förslag på bakåtsteg nekat
takebackPropositionAccepted=Förslag på bakåtsteg godkännt
takebackPropositionCanceled=Förslag på bakåtsteg avbrutet
yourOpponentProposesATakeback=Din motståndare vill ta tillbaka ett drag
bookmarkThisGame=Bokmärk detta spel
toggleBackground=Ställa in bakgrundsfärg
search=Sök
advancedSearch=Avancerad Sökning
tournament=Turnering
tournaments=Turneringar
tournamentPoints=Turneringpoäng
viewTournament=Visa turnering
freeOnlineChessGamePlayChessNowInACleanInterfaceNoRegistrationNoAdsNoPluginRequiredPlayChessWithComputerFriendsOrRandomOpponents=Gratis Schack på internet. Spela Schack nu, med ett enkelt gränssnitt. Ingen registrering, inga annonser, inga instickningsprogram behövs. Spela Schack mot datorn, vänner eller vem som helst.
teams=Lag
nbMembers=%s medlemmar
allTeams=Alla lag
newTeam=Nytt lag
myTeams=Mina lag
noTeamFound=Inget lag funnet
joinTeam=Gå med lag
quitTeam=Lämna lag
anyoneCanJoin=Vem som helst kan gå med
aConfirmationIsRequiredToJoin=Bekräftelse nödvändig för anslutning
joiningPolicy=Anslutningspolicy
teamLeader=Lagledare
teamBestPlayers=Lag bästa spelare
teamRecentMembers=Lag senaste spelare
xJoinedTeamY=%s gick med i lag %s
xCreatedTeamY=%s skapade lag %s
averageElo=Medeltal Elo
location=Plats
settings=Inställningra
filterGames=Filtrera partier
reset=Ställ tillbaka
apply=Använd
leaderboard=Rankinglista
pasteTheFenStringHere=Klistra in FEN-strängen här
pasteThePgnStringHere=Klistra in PGN-koden här
fromPosition=Från position
continueFromHere=Fortsätt härifrån
importGame=Importera parti
nbImportedGames=%s Importerade partier
thisIsAChessCaptcha=Detta är ett schack-CAPTCHA
clickOnTheBoardToMakeYourMove=Bevisa att du är en människa genom att klicka på brädet för att göra ditt drag.
notACheckmate=Inte schackmatt
colorPlaysCheckmateInOne=%s tur; Schackmatt i ett drag
retry=Försök igen
reconnecting=Återansluter
onlineFriends=Vänner online
noFriendsOnline=Inga vänner online
findFriends=Hitta vänner
favoriteOpponents=Favoritmotståndare
follow=Följ
following=Följer
unfollow=Sluta följa
block=Blockera
blocked=Blockerad
unblock=Avblockera
followsYou=Följer dig
xStartedFollowingY=%s började följa %s
nbFollowers=%s följare
nbFollowing=%s följer
more=Mer
memberSince=Medlem sedan
lastLogin=Senast inloggad
challengeToPlay=Utmaning att spela
player=Spelare
list=Lista
graph=Graf
all=Allt
lessThanNbMinutes=Mindre än %s minuter
xToYMinutes=%s till %s minuter
textIsTooShort=Texten är för kort.
textIsTooLong=Texten är för lång.
required=Nödvändig.
addToChrome=Lägg till Chrome
openTournaments=Öppen turneringar
duration=Varaktighet
winner=Vinnare
standing=Ställning
createANewTournament=Skapa en ny turnering
join=Anslut
withdraw=Ge upp
points=Poäng
wins=Vinster
losses=Förluster
winStreak=Vinst serie
createdBy=Skapad av
waitingForNbPlayers=Väntar på %s players
tournamentIsStarting=Turneringen startar
nbMinutesPerSidePlusNbSecondsPerMove=%s minuter/sida + %s sekunder/drag
membersOnly=Endast medlemmar
boardEditor=Brädeditor
startPosition=Starta position
clearBoard=Rensa bord
savePosition=Spara position
loadPosition=Ladda ställning
isPrivate=Privat
reportXToModerators=Rapportera %s till moderatorerna
profile=Profil
editProfile=Ändra profil
firstName=Tilltalsnamn
lastName=Efternamn
biography=Biografi
country=Land
preferences=Inställningar
watchLichessTV=Titta på Lichess TV
previouslyOnLichessTV=Föregående Lichess TV
todaysLeaders=Dagens ledare
onlinePlayers=Spelare online
progressToday=Utveckling i dag
progressThisWeek=Utveckling denna vecka
progressThisMonth=Utveckling denna vecka
leaderboardThisWeek=Utveckling denna vecka
leaderboardThisMonth=Utveckling denna vecka
activeToday=Aktiva i dag
activeThisWeek=Aktiva denna vecka
activePlayers=Aktiva spelare
bestBulletPlayers=Bästa bullet spelare
bestBlitzPlayers=Bästa blitz spelare
bestSlowPlayers=Bästa långsamma spelare
bewareTheGameIsRatedButHasNoClock=OBS! Spelet är rankat men har ingen tidsgräns.
