playWithAFriend=Spela med en vän
inviteAFriendToPlayWithYou=Bjud in en vän att spela med dig
playWithTheMachine=Spela mot datorn
challengeTheArtificialIntelligence=Utmana den artificella intelligensen
toInviteSomeoneToPlayGiveThisUrl=För att bjuda in någon att spela, ge dem den här länken
gameOver=Partiet är slut
waitingForOpponent=Väntar på motståndare
waiting=Väntar
yourTurn=Din tur
aiNameLevelAiLevel=%s nivå %s
level=Nivå
toggleTheChat=Dölj/visa chattrutan
toggleSound=Ljud av/på
chat=Chatt
resign=Ge upp
checkmate=Schackmatt
stalemate=Stallmatt
white=Vit
black=Svart
createAGame=Skapa ett parti
noGameAvailableRightNowCreateOne=Inget spel tillgängligt just nu, skapa ett!
whiteIsVictorious=Vit vinner
blackIsVictorious=Svart vinner
playWithTheSameOpponentAgain=Spela mot samma motståndare igen
newOpponent=Ny moståndare
playWithAnotherOpponent=Spela mot en annan motståndare
yourOpponentWantsToPlayANewGameWithYou=Din motståndare vill spela ett nytt parti med dig
joinTheGame=Anslut till partiet
whitePlays=Vits drag
blackPlays=Svart drag
theOtherPlayerHasLeftTheGameYouCanForceResignationOrWaitForHim=Den andre spelaren har lämnat partiet. Du kan tvinga fram att han ger upp, eller vänta på honom.
makeYourOpponentResign=Tvinga din motståndare att ge upp
forceResignation=Tvinga att ge upp
talkInChat=Prata i chatten
theFirstPersonToComeOnThisUrlWillPlayWithYou=Den första som använder den här länken kommer att spela med dig
whiteCreatesTheGame=Vit startar ett parti
blackCreatesTheGame=Svart startar ett parti
whiteJoinsTheGame=Vit ansluter till partiet
blackJoinsTheGame=Svart ansluter till partiet
whiteResigned=Vit har gett upp
blackResigned=Svart har gett upp
whiteLeftTheGame=Vit har lämnat partiet
blackLeftTheGame=Svart har lämnat partiet
shareThisUrlToLetSpectatorsSeeTheGame=Dela med den här länken så åskådare kan se spelet
youAreViewingThisGameAsASpectator=Du tittar på spelet som åskådare
replayAndAnalyse=Visa repris och analysera
viewGameStats=Visa statistik
flipBoard=Vänd brädet
threefoldRepetition=Trefaldig upprepning
claimADraw=Hävda remi
offerDraw=Föreslå remi
draw=Remi
nbConnectedPlayers=%s anslutna spelare
talkAboutChessAndDiscussLichessFeaturesInTheForum=Snacka om schack och diskutera sidans funktioner i forumet
seeTheGamesBeingPlayedInRealTime=Se de partier som spelas i realtid
gamesBeingPlayedRightNow=Partier som spelas just nu
viewAllNbGames=Visa alla %s partier
viewNbCheckmates=Visa %s  schackmatt
nbBookmarks=%s Bokmärken
nbPopularGames=%s Populära Spel
nbAnalysedGames=%s Spelen Analyserades
bookmarkedByNbPlayers=Bokmärkt av %s spelare
viewInFullSize=Visa i full storlek
logOut=Logga ut
signIn=Logga in
signUp=Registrera dig
people=Människor
games=Partier
forum=Forum
chessPlayers=Schackspelare
minutesPerSide=Minuter per spelare
variant=Variant
timeControl=Tidskontroll
start=Start
username=Användarnamn
password=Lösenord
haveAnAccount=Har du ett konto?
allYouNeedIsAUsernameAndAPassword=Allt du behöver är ett användarnamn och ett lösenord.
learnMoreAboutLichess=Lär mer om Lichess
rank=Rankning
gamesPlayed=Partier spelade
declineInvitation=Avböj inbjudan
cancel=Avbryt
timeOut=Time out
drawOfferSent=Förslag om oavgjort skickat
drawOfferDeclined=Förslag om oavgjort nekat
drawOfferAccepted=Förslag om oavgjort accepterat
drawOfferCanceled=Förslag om oavgjort avbrutet
yourOpponentOffersADraw=Din motståndare föreslår oavgjort
accept=Acceptera
decline=Avböj
playingRightNow=Spelar nu
abortGame=Avsluta parti
gameAborted=Parti avslutat
standard=Standard
unlimited=Obegränsat
mode=Läge
casual=Casual
rated=Poängsatt
thisGameIsRated=Detta parti spelas om ranking
rematch=Ommatch
rematchOfferSent=Förslag om returmatch skickat
rematchOfferAccepted=Förslag om returmatch accepterat
rematchOfferCanceled=Returmatch anbud avbruten
rematchOfferDeclined=Returmatch anbud avböjt
cancelRematchOffer=Neka ommatch förslag
viewRematch=Visa returmatch
play=Spela
inbox=Inkorg
chatRoom=Chattrum
spectatorRoom=Åskådar rum
composeMessage=Sammanställ meddelande
sentMessages=Sända meddelanden
incrementInSeconds=Ökning i sekunder
freeOnlineChess=Gratis Schack på internet
spectators=Åskådare
nbWins=%s vinster
nbLosses=%s förluster
nbDraws=%s remi
exportGames=Exportera spel
color=Färg
eloRange=Elo mellan
giveNbSeconds=Ge  %s sekunder
searchAPlayer=Sök en spelare
whoIsOnline=Vem är online
allPlayers=Alla spelare
namedPlayers=Namngivna spelare
premoveEnabledClickAnywhereToCancel=Preppdrag är möjliggjord-Klicka var som helst för att avbryta
thisPlayerUsesChessComputerAssistance=Den här spelaren använder schackmotor hjälp
opening=Öppning
takeback=Bakåtsteg
proposeATakeback=Föreslå bakåtsteg
takebackPropositionSent=Förslag på bakåtsteg skickat
takebackPropositionDeclined=Förslag på bakåtsteg nekat
takebackPropositionAccepted=Förslag på bakåtsteg godkännt
takebackPropositionCanceled=Förslag på bakåtsteg avbrutet
yourOpponentProposesATakeback=Din motståndare föreslår ett bakåtsteg
bookmarkThisGame=Bokmärk detta spel
toggleBackground=Ställa in bakgrundsfärg
advancedSearch=Avancerad Sökning
tournament=Turnering
freeOnlineChessGamePlayChessNowInACleanInterfaceNoRegistrationNoAdsNoPluginRequiredPlayChessWithComputerFriendsOrRandomOpponents=Gratis Schack på internet. Spela Schack nu, med ett enkelt gränssnitt. Ingen registrering, inga annonser, inga instickningsprogram behövs. Spela Schack mot datorn, vänner eller vem som helst.
teams=Lag
nbMembers=%s medlemmar
allTeams=Alla lag
newTeam=Nytt lag
myTeams=Mina lag
noTeamFound=Inget lag funnet
joinTeam=Anslut till lag
quitTeam=Lämna lag
anyoneCanJoin=Vem som helst kan ansluta
aConfirmationIsRequiredToJoin=Bekräftelse nödvändig för anslutning
joiningPolicy=Anslutningspolicy
teamLeader=Lagledare
teamBestPlayers=Lag bästa spelare
teamRecentMembers=Lag senaste spelare
averageElo=Medeltal ELO
location=Plats
settings=Inställningra
filterGames=Filtrera partier
reset=Ställ tillbaka
apply=Använd
