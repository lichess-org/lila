playWithAFriend=Spela med en vän
playWithTheMachine=Spela mot datorn
toInviteSomeoneToPlayGiveThisUrl=För att bjuda in någon att spela, ge dem den här länken
gameOver=Partiet är slut
waitingForOpponent=Väntar på motståndare
waiting=Väntar
yourTurn=Din tur
aiNameLevelAiLevel=%s nivå %s
level=Nivå
toggleTheChat=Dölj/visa chattrutan
toggleSound=Ljud av/på
chat=Chatt
resign=Ge upp
checkmate=Schackmatt
stalemate=Patt
white=Vit
black=Svart
randomColor=Slumpvis färg
createAGame=Skapa ett parti
whiteIsVictorious=Vit har vunnit
blackIsVictorious=Svart har vunnit
kingInTheCenter=Kungen är i centrum
threeChecks=Tre schackar
raceFinished=Lopp slut
variantEnding=Variantbaserat slut
newOpponent=Ny motståndare
yourOpponentWantsToPlayANewGameWithYou=Din motståndare vill spela ett nytt parti med dig
joinTheGame=Starta partiet
whitePlays=Vits drag
blackPlays=Svarts drag
theOtherPlayerHasLeftTheGameYouCanForceResignationOrWaitForHim=Motståndaren har kanske lämnat partiet. Du kan nu begära vinst, remi eller invänta att motståndaren kommer tillbaka.
makeYourOpponentResign=Tvinga din motståndare att ge upp partiet
forceResignation=Begär vinst
forceDraw=Begär remi
talkInChat=Chatta
theFirstPersonToComeOnThisUrlWillPlayWithYou=Den första som använder den här länken kommer att spela med dig
whiteResigned=Vit har gett upp
blackResigned=Svart har gett upp
whiteLeftTheGame=Vitspelaren har lämnat partiet
blackLeftTheGame=Svartspelaren har lämnat partiet
shareThisUrlToLetSpectatorsSeeTheGame=Dela den här länken till åskådare som vill se partiet
theComputerAnalysisHasFailed=Datoranalysen misslyckades
viewTheComputerAnalysis=Visa datoranalysen
requestAComputerAnalysis=Begär en datoranalys
computerAnalysis=Datoranalys
analysis=Analys
blunders=Blundrar
mistakes=Misstag
inaccuracies=Felaktigheter
moveTimes=Dragtider
flipBoard=Vänd brädet
threefoldRepetition=Trefaldig repetition
claimADraw=Begär remi
offerDraw=Föreslå remi
draw=Remi
nbConnectedPlayers=%s spelare
gamesBeingPlayedRightNow=Pågående partier
viewAllNbGames=%s partier
viewNbCheckmates=Visa %s schackmatt
nbBookmarks=%s Bokmärken
nbPopularGames=%s Populära partier
nbAnalysedGames=%s Analyserade partier
bookmarkedByNbPlayers=Bokmärkt av %s spelare
viewInFullSize=Visa i full storlek
logOut=Logga ut
signIn=Logga in
newToLichess=Ny användare?
youNeedAnAccountToDoThat=Du behöver ett konto för att göra detta
signUp=Registrera dig
computersAreNotAllowedToPlay=Datorer och datorhjälp är inte tillåtet att spela med. Vänligen, ta inte hjälp ifrån schackmotorer, databaser eller från andra spelare när du spelar. Notera även att skapande av flera konton avskräcks och överdrivet skapande leder till avstängning.
games=Partier
forum=Forum
xPostedInForumY=%s postade i forumet %s
latestForumPosts=Senaste foruminläggen
players=Spelare
minutesPerSide=Minuter per spelare
variant=Variant
variants=Varianter
timeControl=Tidskontroll
realTime=Realtid
correspondence=Korrespondens
daysPerTurn=Dagar per drag
oneDay=En dag
nbDays=%s dagar
nbHours=%s timmar
time=Tid
rating=Rating
ratingStats=Rating statistik
username=Användar namn
usernameOrEmail=Användarnamn
password=Lösenord
haveAnAccount=Har du ett konto?
changePassword=Ändra lösenord
changeEmail=Ändra E-post
email=E-post
emailIsOptional=E-post är valfritt. Lichess kan använda den för att återställa ditt lösenord om du glömmer det.
passwordReset=Återställ lösenord
forgotPassword=Glömt lösenord?
rank=Rankning
gamesPlayed=Partier spelade
nbGamesWithYou=%s partier med dig
declineInvitation=Avböj inbjudan
cancel=Avbryt
timeOut=Tidsförlust
drawOfferSent=Remierbjudande skickat
drawOfferDeclined=Remi avböjd
drawOfferAccepted=Remi accepterad
drawOfferCanceled=Remiförfrågan avbruten
whiteOffersDraw=Vit erbjuder remi
blackOffersDraw=Svart erbjuder remi
whiteDeclinesDraw=Vit avböjer remi
blackDeclinesDraw=Svart avböjer remi
yourOpponentOffersADraw=Din motståndare erbjuder remi
accept=Acceptera
decline=Avböj
playingRightNow=Spelar parti just nu
finished=Avslutade
abortGame=Avbryt partiet
gameAborted=Partiet avbröts
standard=Standard
unlimited=Obegränsad
mode=Läge
casual=Ej rankat
rated=Rankat
thisGameIsRated=Detta parti är rankat
rematch=Returmatch
rematchOfferSent=Förslag om returmatch skickat
rematchOfferAccepted=Förslag om returmatch accepterat
rematchOfferCanceled=Anbud om returmatch upphävt
rematchOfferDeclined=Anbud om returmatch avböjt
cancelRematchOffer=Upphäv returmatchförslag
viewRematch=Visa returmatch
play=Spela
inbox=Inkorg
chatRoom=Chattrum
spectatorRoom=Åskådarrum
composeMessage=Skriv meddelande
noNewMessages=Inga nya meddelanden
subject=Ämne
recipient=Mottagare
send=Skicka
incrementInSeconds=Tilläggssekunder
freeOnlineChess=Gratis schack på internet
spectators=Åskådare
nbWins=%s vinster
nbLosses=%s förluster
nbDraws=%s remier
exportGames=Exportera spel
ratingRange=Ratingomfång
giveNbSeconds=Ge  %s sekunder
premoveEnabledClickAnywhereToCancel=Premove aktiverat - Klicka var som helst för att avbryta
thisPlayerUsesChessComputerAssistance=Den här spelaren tar hjälp av schackmotor
thisPlayerArtificiallyIncreasesTheirRating=Den här spelaren ökar/minskar sin rating artificiellt
opening=Öppning
openingExplorer=Åbning opdagelse
takeback=Gör om drag
proposeATakeback=Frågar motståndaren om du får göra om draget
takebackPropositionSent=Förslag att göra om draget skickat
takebackPropositionDeclined=Förslag att göra om draget nekat av motståndaren
takebackPropositionAccepted=Förslag att göra om draget godkänt
takebackPropositionCanceled=Förslag på att göra om draget har dragits tillbaka
yourOpponentProposesATakeback=Din motståndare vill göra om det senaste draget
bookmarkThisGame=Bokmärk detta parti
search=Sök
advancedSearch=Avancerad sökning
tournament=Turnering
tournaments=Turneringar
tournamentPoints=Turneringspoäng
viewTournament=Visa turnering
backToTournament=Tillbaka till turnering
backToGame=Tillbaka till partiet
freeOnlineChessGamePlayChessNowInACleanInterfaceNoRegistrationNoAdsNoPluginRequiredPlayChessWithComputerFriendsOrRandomOpponents=Gratis Schack på internet. Spela Schack nu, med ett enkelt gränssnitt. Ingen registrering, inga annonser, inga instickningsprogram behövs. Spela Schack mot datorn, vänner eller vem som helst.
teams=Lag
nbMembers=%s medlemmar
allTeams=Alla lag
newTeam=Nytt lag
myTeams=Mina lag
noTeamFound=Inget lag hittat
joinTeam=Gå med i lag
quitTeam=Lämna lag
anyoneCanJoin=Vem som helst kan gå med
aConfirmationIsRequiredToJoin=Bekräftelse nödvändig för att gå med
joiningPolicy=Deltagningspolicy
teamLeader=Lagledare
teamBestPlayers=Topplista
teamRecentMembers=Nya medlemmar
xJoinedTeamY=%s gick med i lag %s
xCreatedTeamY=%s skapade lag %s
averageElo=Medelrating
location=Plats
settings=Inställningar
filterGames=Filtrera partier
reset=Återställ
apply=Använd
leaderboard=Rankinglista
pasteTheFenStringHere=Klistra in FEN-koden här
pasteThePgnStringHere=Klistra in PGN-koden här
fromPosition=Från position
continueFromHere=Fortsätt härifrån
importGame=Importera parti
nbImportedGames=%s Importerade partier
thisIsAChessCaptcha=Detta är en schack-CAPTCHA
clickOnTheBoardToMakeYourMove=Bevisa att du är en människa genom att klicka på brädet och göra ditt drag.
notACheckmate=Inte schackmatt
colorPlaysCheckmateInOne=%s tur; Schackmatt i ett drag
retry=Försök igen
reconnecting=Återansluter
onlineFriends=Vänner online
noFriendsOnline=Inga vänner online
findFriends=Hitta vänner
favoriteOpponents=Favoritmotståndare
follow=Följ
following=Följer
unfollow=Sluta följa
block=Blockera
blocked=Blockerad
unblock=Avblockera
followsYou=Följer dig
xStartedFollowingY=%s började följa %s
nbFollowers=%s följare
nbFollowing=%s följer
more=Mer
memberSince=Medlem sedan
lastLogin=Senast inloggad
challengeToPlay=Utmana till ett spel
player=Spelare
list=Lista
graph=Graf
lessThanNbMinutes=Mindre än %s minuter
xToYMinutes=%s till %s minuter
textIsTooShort=Texten är för kort.
textIsTooLong=Texten är för lång.
required=Obligatoriskt.
openTournaments=Öppna turneringar
duration=Varaktighet
winner=Vinnare
standing=Ställning
createANewTournament=Skapa en ny turnering
join=Delta
withdraw=Lämna
points=Poäng
wins=Vinster
losses=Förluster
winStreak=Vinstserie
createdBy=Skapad av
tournamentIsStarting=Turneringen startar
membersOnly=Endast medlemmar
boardEditor=Brädeditor
startPosition=Startposition
clearBoard=Rensa bräde
savePosition=Spara ställning
loadPosition=Ladda ställning
isPrivate=Privat
reportXToModerators=Rapportera %s till moderatorerna
profile=Profil
editProfile=Ändra profil
firstName=Förnamn
lastName=Efternamn
biography=Biografi
country=Land
preferences=Inställningar
watchLichessTV=Titta på Lichess TV
previouslyOnLichessTV=Föregående Lichess TV
onlinePlayers=Spelare online
activeToday=Aktivast i dag
activePlayers=Aktiva spelare
bewareTheGameIsRatedButHasNoClock=OBS! Spelet är rankat men har ingen tidsgräns.
training=Träning
yourPuzzleRatingX=Din problemlösarrating: %s
findTheBestMoveForWhite=Hitta bästa draget för vit.
findTheBestMoveForBlack=Hitta bästa draget för svart.
toTrackYourProgress=För att följa din utveckling:
trainingSignupExplanation=Lichess kommer att erbjuda schackproblem som matchar din förmåga, vilket ger dig bättre träning.
recentlyPlayedPuzzles=Nyligen spelade schackproblem
puzzleId=Schackproblem %s
puzzleOfTheDay=Dagens schackproblem
clickToSolve=Klicka för att lösa
goodMove=Bra drag
butYouCanDoBetter=Men det finns ännu bättre drag.
bestMove=Bästa draget!
keepGoing=Fortsätt...
puzzleFailed=Feldrag
butYouCanKeepTrying=Men du kan fortsätta försöka.
victory=Rätt!
giveUp=Ge upp
puzzleSolvedInXSeconds=Schackproblemet löstes på %s sekunder.
wasThisPuzzleAnyGood=Var det här schackproblemet bra?
pleaseVotePuzzle=Hjälp lichess att bli bättre genom att rösta (använd pil upp eller pil ner):
thankYou=Tack!
ratingX=Rating: %s
playedXTimes=Spelat %s gånger
fromGameLink=Från parti: %s
startTraining=Starta träning
continueTraining=Fortsätt träning
retryThisPuzzle=Testa detta schackproblem igen
thisPuzzleIsCorrect=Det här schackproblemet är korrekt och intressant
thisPuzzleIsWrong=Det här schackproblemet är fel eller tråkigt
youHaveNbSecondsToMakeYourFirstMove=du har %s sekunder för att göra första draget
nbGamesInPlay=%s partier spelas
automaticallyProceedToNextGameAfterMoving=Gör att du automatiskt fortsätter till nästa parti efter du gjort ett drag
autoSwitch=Automatiskt partibyte
openingId=Öppning %s
yourOpeningRatingX=Din öppningsrating: %s
findNbStrongMoves=Hitta %s starka drag
thisMoveGivesYourOpponentTheAdvantage=Detta drag ger din motståndare övertaget
openingFailed=Misslyckad öppning
openingSolved=Öppning löst
recentlyPlayedOpenings=Nyligen spelade öppningar
puzzles=Problemlösningar
coordinates=Koordinater
openings=Öppningar
latestUpdates=Senaste uppdateringarna
tournamentWinners=Turneringsvinnare
name=Namn
description=Beskrivning
no=Nej
yes=Ja
help=Hjälp:
createANewTopic=Skapa ett nytt ämne
topics=Ämnen
posts=Inlägg
lastPost=Senaste inlägget
views=Visningar
replies=Svar
replyToThisTopic=Svara på ämnet
reply=Svara
message=Meddelande
createTheTopic=Skapa ämnet
reportAUser=Rapportera en användare
user=Användare
reason=Anledning
whatIsIheMatter=Vad är problemet?
cheat=Fusk
insult=Förolämpning
troll=Troll
other=Övrigt
reportDescriptionHelp=Klistra in länken till spelet och förklara vad som är fel med den här användarens beteende.
by=av %s
thisTopicIsNowClosed=Det här ämnet är nu stängt.
theming=Teman
donate=Donera
blog=Blogg
questionsAndAnswers=Frågor & Svar
notes=Anteckningar
typePrivateNotesHere=Skriv privata anteckningar här
gameDisplay=Spelutseende
pieceAnimation=Pjäsanimation
materialDifference=Materialskillnad
closeAccount=Avsluta konto
closeYourAccount=Avsluta ditt konto
changedMindDoNotCloseAccount=Jag ändrade mig, avsluta inte mitt konto
closeAccountExplanation=Är du säker att du vill avsluta ditt konto? Att avsluta ditt konto är ett permanent beslut. Du kommer inte längre kunna logga in och din profilsida kommer inte längre vara tillgänglig.
thisAccountIsClosed=Det här kontot är avslutat
invalidUsernameOrPassword=Ogiltigt användarnamn eller lösenord
emailMeALink=Maila mig en länk
currentPassword=Nuvarande lösenord
newPassword=Nytt lösenord
newPasswordAgain=Repetera lösenord
boardHighlights=Brädmarkeringar (föregående drag och schack)
pieceDestinations=Möjliga drag (giltiga drag och premoves)
boardCoordinates=Brädkoordinater (A-H, 1-8)
moveListWhilePlaying=Lista med drag under spelets gång
chessClock=Schack-klocka
tenthsOfSeconds=Tiondels sekunder
never=Aldrig
whenTimeRemainingLessThanTenSeconds=När återstående tid < 10 sekunder
horizontalGreenProgressBars=Horisontella gröna förloppsindikatorer
soundWhenTimeGetsCritical=Ljud när tiden blir kritisk
gameBehavior=Spelbeteende
premovesPlayingDuringOpponentTurn=Premoves (göra drag i förväg under motståndarens tur)
takebacksWithOpponentApproval=Ta tillbaka drag (med motståndarens godkännande)
promoteToQueenAutomatically=Uppgradera till drottning automatiskt
claimDrawOnThreefoldRepetitionAutomatically=Begär oavgjort automatiskt vid %strefaldig upprepning%s
privacy=Sekretess
letOtherPlayersFollowYou=Låt andra spelare följa dig
letOtherPlayersChallengeYou=Låt andra spelare utmana dig
sound=Ljud
soundControlInTheTopBarOfEveryPage=Ljudkontrollen finns längst till höger i den översta menyn på varje sida.
yourPreferencesHaveBeenSaved=Dina inställningar har sparats.
none=Ingen
fast=Snabb
normal=Medel
slow=Långsam
insideTheBoard=På brädet
outsideTheBoard=Utanför brädet
onSlowGames=På långsamma spel
always=Alltid
inCasualGamesOnly=Endast i icke rankade spel
whenPremoving=Vid premove
whenTimeRemainingLessThanThirtySeconds=När återstående tid < 30 sekunder
difficultyEasy=Lätt
difficultyNormal=Medel
difficultyHard=Svår
xLeftANoteOnY=%s skrev en notering på %s
xCompetesInY=%s tävlar i %s
xAskedY=%s frågade %s
xAnsweredY=%s svarade %s
xCommentedY=%s kommenterade %s
timeline=Tidslinje
seeAllTournaments=Se alla turneringar
starting=Startar:
allInformationIsPublicAndOptional=All information är allmän och frivillig.
yourCityRegionOrDepartment=Din stad, region eller område.
biographyDescription=Berätta om dig själv, vad du gillar med schack, dina favoritöppningar, spel, spelare…
maximumNbCharacters=Max: %s tecken.
blocks=%s blockeringar
listBlockedPlayers=Lista spelare som du blockerat
human=Människa
computer=Dator
side=Sida
clock=Klocka
unauthorizedError=Tillgång är oauktoriserad
noInternetConnection=Ingen internet förbindelse. Du kan spela offline från menyn
connectedToLichess=Du är nu ansluten till lichess.org
signedOut=Du har loggat ut
loginSuccessful=Lyckad inloggning
playOnTheBoardOffline=Spela offline, över bräden
playOfflineComputer=Spela mot dator offline
opponent=Motståndare
learn=Lära sig
community=Gemenskap
tools=Verktyg
increment=Tillägg
board=Bräde
pieces=Pjäser
sharePGN=Dela PGN
playOnline=Spela online
playOffline=Spela offline
allowAnalytics=Tillåt anonym statistik
shareGameURL=Dela parti-URL
error.required=Detta fältet är obligatoriskt
error.email=Ogiltig e-postadress
error.email_acceptable=Oacceptabel e-postadress
error.email_unique=Det finns redan ett konto med denna e-postadress
blindfoldChess=Blindschack (Osynliga pjäser)
moveConfirmation=Bekräftelse av drag
inCorrespondenceGames=I korrespondensparti
ifRatingIsPlusMinusX=Om rating är ± %s
onlyFriends=Bara vänner
menu=Meny
castling=Rockad
whiteCastlingKingside=Vit O-O
whiteCastlingQueenside=Vit O-O-O
blackCastlingKingside=Svart O-O
blackCastlingQueenside=Svart O-O-O
nbForumPosts=%s av foruminlägg
tpTimeSpentPlaying=Total speltid: %s
watchGames=Titta på spel
tpTimeSpentOnTV=Total TV-tid: %s
watch=Titta
internationalEvents=Internationella evenemang
videoLibrary=Videobibliotek
mobileApp=Mobilapp
webmasters=Webbmasters
contribute=Hjälp till
contact=Kontakt
termsOfService=Användarvillkor
sourceCode=Källkod
simultaneousExhibitions=Simultanschack
host=Värd
createdSimuls=Nyligen skapade simuls
hostANewSimul=Skapa ny simul
noSimulFound=Simul hittades ej
noSimulExplanation=Denna simul existerar inte.
returnToSimulHomepage=Återvänd till hemsidan för simul
aboutSimul=Simuls går ut på att en spelare möter flera spelare samtidigt.
aboutSimulImage=Av totalt 50 partier vann Fischer 47, spelade lika två och förlorade en.
aboutSimulRealLife=Konceptet är taget från verkliga evenemang. I verkligheten involverar det att simul-värden rör sig från bord till bord för att göra sina drag.
aboutSimulRules=När simultanen börjar startar varje spelare ett parti med värden som spelar vit i alla partier.  Simultanen slutar när alla partier är avklarade.
aboutSimulSettings=Simultanpartier är alltid orankade. Returmatch, ångerdrag och "extratid" är inaktiverat.
create=Skapa
whenCreateSimul=När du skapar en simul får du spela mot flera spelare samtidigt.
simulVariantsHint=Om du väljer flera varianter får varje spelare välja vilken de vill spela.
simulClockHint=Inställningar för fischerklocka. Ju fler spelare du tar dig an, desto mer tid kan du behöva.
simulAddExtraTime=Du kan lägga till extra tid för att klara av simultanspelet.
simulHostExtraTime=Värdens extratid
lichessTournaments=Lichess-turneringar
tournamentFAQ=Turnering FAQ
tournamentOfficial=Officiell
timeBeforeTournamentStarts=Tid tills turneringen börjar
averageCentipawnLoss=Genomsnittligt förlorad hundradelsbonde
keyboardShortcuts=Snabbkommandon
keyMoveBackwardOrForward=bakåtdrag/framåtdrag
keyGoToStartOrEnd=gå till början/slut
keyShowOrHideComments=Visa/göm kommentarer
keyEnterOrExitVariation=påbörja/avsluta variant
keyYouCanDrawArrowsCirclesAndScrollToMove=Tryck ned shift och klicka (alternativt högerklicka) för att rita ut cirklar eller pilar på brädet. Du kan också skrolla över brädet för att göra drag i partiet.
newTournament=Ny turnering
tournamentHomeTitle=Schackturnering med olika betänketider och schackvarianter
tournamentHomeDescription=Spela snabba schackturneringar! Delta i en officiell planerad turnering, eller skapa din egen. Bullet, Blitz, Classical, Chess960, King of the Hill, Threecheck och fler alternativ erbjuds för ändlöst schackskoj.
tournamentNotFound=Turnering ej funnen
tournamentDoesNotExist=Denna turnering finns inte
tournamentMayHaveBeenCanceled=Den kan ha blivit inställd om alla spelare lämnade den innan start.
returnToTournamentsHomepage=Återgå till turneringens hemsida
weeklyPerfTypeRatingDistribution=Månatlig %s rating fördelning
nbPerfTypePlayersThisWeek=%s %s spelare denna månad.
yourPerfTypeRatingisRating=Din %s rating är %s.
youAreBetterThanPercentOfPerfTypePlayers=Du är bättre än %s av %s spelarna.
youDoNotHaveAnEstablishedPerfTypeRating=Du har inte en etablerad %s rating.
checkYourEmail=Kolla din email
weHaveSentYouAnEmailClickTheLink=Vi har skickat ett e-postmeddelande . Klicka på länken i meddelandet för att aktivera ditt konto.
ifYouDoNotSeeTheEmailCheckOtherPlaces=Om du inte ser e-post, kontrollera andra ställen kan det vara, som ditt skräp, spam, sociala eller andra mappar.
areYouSureYouEvenRegisteredYourEmailOnLichess=Är du säker på att du även registrerat din e-post på lichess?
itWasNotRequiredForYourRegistration=Det var inte obligatorisk/ett krav för din registrering
weHaveSentYouAnEmailTo=Vi har skickat ett e-postmeddelande till %s.Tryck på länken i eposten för att återställa ditt lösenord.
byRegisteringYouAgreeToBeBoundByOur=Genom att registrera samtycker du till att vara bunden av våra %s.
networkLagBetweenYouAndLichess=Nätverks fördröjning mellan dig och lichess
timeToProcessAMoveOnLichessServer=Tid att bearbeta ett drag på lichess server
downloadAnnotated=nedladdning kommenterad
downloadRaw=Hämta rå
downloadImported=nedladdning importeras
printFriendlyPDF=Utskriftsvänlig PDF
crosstable=tvär Tabell
youCanAlsoScrollOverTheBoardToMoveInTheGame=Du kan också rulla över styrelsen att röra sig i spelet.
pressShiftPlusClickOrRightClickToDrawCirclesAndArrowsOnTheBoard=Tryck på Skift + klicka eller högerklicka för att rita cirklar och pilar på tavlan.
confirmResignation=Bekräfta resignation
letOtherPlayersMessageYou=Tillåt andra spelare att skicka meddelanden till dig
shareYourInsightsData=Dela din inblicksinformation
youHaveAlreadyRegisteredTheEmail=Du har redan registrerat en email adress: %s
kidMode=Barnsäkert läge
playChessEverywhere=Spela schack överallt
asFreeAsLichess=Lika gratis som lichess
builtForTheLoveOfChessNotMoney=Skapad med kärlek för schack, inte pengar
zeroAdvertisement=Ingen reklam
phoneAndTablet=Mobil och surfplatta
correspondenceChess=Korrespondensschack
